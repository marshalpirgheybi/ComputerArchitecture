module
    
    endmodule