module
    
endmodule