module a (in,out);
    input a;
    output out;
endmodule